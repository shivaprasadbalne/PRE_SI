module ASYNC_FIFO#(parameter FIFO_DEPTH = 8,)(
input DATA_IN, 
input WRITE_EN, 
input WRITE_PTR, 
input WRITE_CLK;
output

);